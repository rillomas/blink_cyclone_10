module FullAdder(
	input logic a,
	input logic b,
	input logic ci,
	output logic s,
	output logic co);
	logic s0, co0, co1;
	HalfAdder ha_before(.a(a), .b(b), .s(s0), .co(co0));
	HalfAdder ha_after(.a(s0), .b(ci), .s(s), .co(co1));
	assign co = co0 | co1;
endmodule